LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
ENTITY T_FF_tb IS
END T_FF_tb;
 
ARCHITECTURE behavior OF T_FF_tb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT T_FF
    PORT(
         T_input : IN  std_logic;
         clk : IN  std_logic;
         rst : IN  std_logic;
         T_output : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal T_input : std_logic := '1';
   signal clk : std_logic := '0';
   signal rst : std_logic := '1';

 	--Outputs
   signal T_output : std_logic;

   -- Clock period definitions
   constant clk_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: T_FF PORT MAP (
          T_input => T_input,
          clk => clk,
          rst => rst,
          T_output => T_output
        );

   -- Clock process definitions
   clk_process :process
   begin
		clk <= '0';
		wait for clk_period/2;
		clk <= '1';
		wait for clk_period/2;
   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      wait for clk_period*10;
		
		rst <= '0';
		wait for 10 ns;
    
		
      T_input <= '0';
		wait for 10 ns;
		
      T_input <= '1';
		wait for 60 ns;
		
		rst <= '1';

      wait;
   end process;

END;

