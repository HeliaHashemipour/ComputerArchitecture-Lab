------------------------------
--Lab04-Ripple Carry Adder
------------------------------
library ieee;
use ieee.std_logic_1164.all;

 Entity half_adder IS
 Port(
	A: IN std_logic;
	B: IN std_logic;
	S: OUT std_logic;
	Cout : OUT std_logic);
 End Entity half_adder;

 Architecture Behavioral of half_adder IS
begin
	S <= A xor B;
	Cout <= A and B;
	
end Behavioral;
